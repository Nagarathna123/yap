//Control unit

//macros
//instruction width
`define INSTRUCTION_WIDTH 32
//ALU control signal width
`define ALU_CTRL_WIDTH 5

//Instruction types
//R-type
`define R_TYPE 5'b01100
//I-type
`define JALR 5'b11001
`define LOAD 5'b00000
`define ALU 5'b00100
//S-type
`define STORE 5'b01000
//SB-type
`define BRANCH 5'b11000
//U-type
`define U_TYPE 5'b01101, 5'b00101
//UJ-type
`define JAL 5'b11011

module ctrl(
	//outputs
	/*ALU control signal
	bits 2 - 0 : ALU operation to be performed
	bit 3 : Set to 1 when a subtract operation is to be performed
	bit 4 : Set to 1 in case of branch instruction
	*/
	output reg [(`ALU_CTRL_WIDTH-1):0] alu_ctrl,
	//Register file write enable signal
	output reg reg_file_wr_en,
	/*Register file writeback select signal (2 bits)
	(00) output of ALU
	(01) output of data memory
	(10) output of PC+4
	(11) output of PC+immediate value
	*/
	output reg [1:0] reg_file_wr_back_sel,
	//ALU operand select signal
	output reg alu_op2_sel,
	//Data memory read enable signal
	output reg d_mem_rd_en,
	//Data memory write enalbe signal
	output reg d_mem_wr_en,
	/*Data memory size
	(00) 32 bit value
	(01) 16 bit value
	(10) 8 bit value
	(11) undefined
	*/
	output reg [2:0] d_mem_size,
	//JAL instruction
	output reg jal,
	//JALR instruction
	output reg jalr, 
	//inputs
	input [(`INSTRUCTION_WIDTH - 1):0] inst
);
	
	//combinational logic
	always @ (*) begin
		//first check if the input instruction is valid
		if (inst[1:0] == 2'b11) begin
			//determine the type of instruction
			case (inst[6:2])
			
				//R-type
				`R_TYPE: begin
					//set the alu_ctrl signal to be the packed version of
					//MSB = inst[31] and remaining bits = funct3 field as specified in the ISA
					//MSB = 1 distinguishes between SUB and ADD
					//MSB = 1 ==> SUB
					//ALU control signal
					alu_ctrl[3:0] = {inst[30], inst[14:12]};
					//no branching
					alu_ctrl[4] = 1'b0;
					//Register file write enable signal
					//the value generated from the ALU is always written back to the register file in R-type
					reg_file_wr_en = 1'b1;
					//Register file writeback select signal
					//by default, the value generated by the ALU is written back 
					reg_file_wr_back_sel = 2'b00;
					//ALU operand select signal
					//the second operand for the ALU is obtained from the register file
					alu_op2_sel = 1'b0;
					//Data memory read enable signal
					//Data memory is not read
					data_mem_rd_en = 1'b0;
					//Data memory write enalbe signal
					//Data memory is not written to
					data_mem_wr_en = 1'b0;
					//No data is written to data memory
					//set to default value
					d_mem_size = 2'b00;
					//JAL instruction
					//not valid
					jal = 1'b0;
					//JALR instruction
					//not valid
					jalr = 1'b0;
				end
				
				//I-type
				`LOAD: begin
					//ALU control signal
					//set the ALU control to add operation
					//The operand obtained from the register is added to the immediate value
					//no branching
					alu_ctrl = {(`ALU_CTRL_WIDTH){1'b0}};
					//Register file write enable signal
					//Value read from the data memory is written back to the register file
					reg_file_wr_en = 1'b1;
					//Register file writeback select signal
					//Value read from data memory is written back to register file
					reg_file_wr_back_sel = 2'b01;
					//ALU operand select signal
					//select the sign or zero extended operand
					alu_op2_sel = 1'b1;
					//Data memory read enable signal
					//The value is loaded from data memory
					data_mem_rd_en = 1'b1;
					//Data memory write enalbe signal
					//no value is written to data memory
					data_mem_wr_en = 1'b0;
					//data is written to data memory
					//size depends on 
					d_mem_size = 2'b00;
					//JAL instruction
					//not valid
					jal = 1'b0;
					//JALR instruction
					//not valid
					jalr = 1'b0;
				end
				
				`ALU: begin
					//ALU control signal
					//set the alu_ctrl signal to {1'b0, "funct3"}
					//MSB = 1'b0, no subtract instructions
					alu_ctrl = {1'b0, inst[14:12]};
					//Register file write enable signal
					//value generated by the ALU is always written back to the register file
					reg_file_wr_en = 1'b1;
					//Register file writeback select signal
					//select the value generated by the ALU
					reg_file_wr_back_sel = 1'b0;
					//ALU operand select signal
					//select the sign or zero extended immediate value
					alu_op2_sel = 1'b1;
					//Data memory read enable signal
					//no value is read from data memory
					data_mem_rd_en = 1'b0;
					//Data memory write enalbe signal
					//no value is written back to data memory
					data_mem_wr_en = 1'b0;	
				end	
				
				//S-type
				`STORE: begin
					//ALU control signal
					//set the ALU control signal to add "rs1" to immediate value
					alu_ctrl = {(`ALU_CTRL_WIDTH){1'b0}};
					//Register file write enable signal
					//no write to register file
					reg_file_wr_en = 1'b0;
					//Register file writeback select signal
					//signal value does not matter
					reg_file_wr_back_sel = 1'b0;
					//ALU operand select signal
					//select the sign or zero extended immediate value
					alu_op2_sel = 1'b1;
					//Data memory read enable signal
					//no data is read from data memory
					data_mem_rd_en = 1'b0;
					//Data memory write enalbe signal
					//Data is written to data memory
					data_mem_wr_en = 1'b1;
				end
				
				//default
				default: begin
					//set all signals to default value (0)
					//ALU control signal
					alu_ctrl = {(`ALU_CTRL_WIDTH){1'b0}};
					//Register file write enable signal
					reg_file_wr_en = 1'b0;
					//Register file writeback select signal
					reg_file_wr_back_sel = 1'b0;
					//ALU operand select signal
					alu_op2_sel = 1'b0;
					//Data memory read enable signal
					data_mem_rd_en = 1'b0;
					//Data memory write enalbe signal
					data_mem_wr_en = 1'b0;
				end
			
			endcase
		end
		
		else begin
			//set all signals to default value (0)
			//ALU control signal
			alu_ctrl = {(`ALU_CTRL_WIDTH){1'b0}};
			//Register file write enable signal
			reg_file_wr_en = 1'b0;
			//Register file writeback select signal
			reg_file_wr_back_sel = 1'b0;
			//ALU operand select signal
			alu_op2_sel = 1'b0;
			//Data memory read enable signal
			data_mem_rd_en = 1'b0;
			//Data memory write enalbe signal
			data_mem_wr_en = 1'b0;
		end
	end

endmodule
